module encrypt(
    output [255:0] ct,
    input [255:0] pt,
    input [63:0] key
);
endmodule

module decrypt(
    output [255:0] ct,
    input [255:0] pt,
    input [63:0] key
);
endmodule

module padd(
    output [255:0] ct,
    input 
);
endmodule

module keygen();
endmodule

module alu64bit();
endmodule

module algotest();
endmodule